LIBRARY ieee;
LIBRARY STD;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
USE STD.textio.all;
USE ieee.std_logic_textio.all;

package helper_funcs is
  subtype static_char is character;
  function char2ascii(char : static_char) return STD_LOGIC_VECTOR;
end helper_funcs;

package body helper_funcs is
  function char2ascii(char : static_char) return STD_LOGIC_VECTOR is
  variable ascii : STD_LOGIC_VECTOR(7 downto 0);
  variable v_char : static_char;
  begin
    v_char  := char;
    case v_char is
      when ' '    => ascii := x"20";
      when 'a'    => ascii := x"61";
      when 'b'    => ascii := x"62";
      when 'c'    => ascii := x"63";
      when 'd'    => ascii := x"64";
      when 'e'    => ascii := x"65";
      when 'f'    => ascii := x"66";
      when 'g'    => ascii := x"67";
      when 'h'    => ascii := x"68";
      when 'i'    => ascii := x"69";
      when 'j'    => ascii := x"6A";
      when 'k'    => ascii := x"6B";
      when 'l'    => ascii := x"6C";
      when 'm'    => ascii := x"6D";
      when 'n'    => ascii := x"6E";
      when 'o'    => ascii := x"6F";
      when 'p'    => ascii := x"70";
      when 'q'    => ascii := x"71";
      when 'r'    => ascii := x"72";
      when 's'    => ascii := x"73";
      when 't'    => ascii := x"74";
      when 'u'    => ascii := x"75";
      when 'v'    => ascii := x"76";
      when 'w'    => ascii := x"77";
      when 'x'    => ascii := x"78";
      when 'y'    => ascii := x"79";
      when 'z'    => ascii := x"7A";
      when 'A'    => ascii := x"41";
      when 'B'    => ascii := x"42";
      when 'C'    => ascii := x"43";
      when 'D'    => ascii := x"44";
      when 'E'    => ascii := x"45";
      when 'F'    => ascii := x"46";
      when 'G'    => ascii := x"47";
      when 'H'    => ascii := x"48";
      when 'I'    => ascii := x"49";
      when 'J'    => ascii := x"4A";
      when 'K'    => ascii := x"4B";
      when 'L'    => ascii := x"4C";
      when 'M'    => ascii := x"4D";
      when 'N'    => ascii := x"4E";
      when 'O'    => ascii := x"4F";
      when 'P'    => ascii := x"50";
      when 'Q'    => ascii := x"51";
      when 'R'    => ascii := x"52";
      when 'S'    => ascii := x"53";
      when 'T'    => ascii := x"54";
      when 'U'    => ascii := x"55";
      when 'V'    => ascii := x"56";
      when 'W'    => ascii := x"57";
      when 'X'    => ascii := x"58";
      when 'Y'    => ascii := x"59";
      when 'Z'    => ascii := x"5A";
      when '!'    => ascii := x"21";
      --when '\"'   => ascii := x"22";
      when '#'    => ascii := x"23";
      when '$'    => ascii := x"24";
      when '%'    => ascii := x"25";
      when '&'    => ascii := x"26";
      when '('    => ascii := x"28";
      when ')'    => ascii := x"29";
      when '*'    => ascii := x"2A";
      when '+'    => ascii := x"2B";
      when ':'    => ascii := x"3A";
      when '<'    => ascii := x"3C";
      when '>'    => ascii := x"3E";
      when '?'    => ascii := x"3F";
      when '@'    => ascii := x"40";
      when '^'    => ascii := x"5E";
      when '_'    => ascii := x"5F";
      when '{'    => ascii := x"7B";
      when '|'    => ascii := x"7C";
      when '}'    => ascii := x"7D";
      when '~'    => ascii := x"7E";
      when '0'    => ascii := x"30";
      when '1'    => ascii := x"31";
      when '2'    => ascii := x"32";
      when '3'    => ascii := x"33";
      when '4'    => ascii := x"34";
      when '5'    => ascii := x"35";
      when '6'    => ascii := x"36";
      when '7'    => ascii := x"37";
      when '8'    => ascii := x"38";
      when '9'    => ascii := x"39";
      when '''    => ascii := x"27";
      when ','    => ascii := x"2C";
      when '-'    => ascii := x"2D";
      when '.'    => ascii := x"2E";
      when '/'    => ascii := x"2F";
      when ';'    => ascii := x"3B";
      when '='    => ascii := x"3D";
      when '['    => ascii := x"5B";
      --when "\"    => ascii := x"5C";
      when ']'    => ascii := x"5D";
      when '`'    => ascii := x"60";
      when others => NULL;
    end case;
    return ascii;
  end function;
end helper_funcs;
